// instruction decode unit

`include "defines.svh"

module decode (
    input  logic [31:0] instr,

    output logic [3:0]  rd,
    output logic [3:0]  rs1,
    output logic [3:0]  rs2,

    output logic        is_alu_op, // TODO drive this
    output alu_op_t     alu_op,
    output comp_t       comp_op,
    output logic        subtract,
    output logic        shift_right,
    output logic        shift_arith,
    output logic        is_auipc,
    
    output logic        is_load_op,
    output load_op_t    load_op,
    output logic        is_store_op,
    output store_op_t   store_op,

    output logic        is_br_type,
    output br_type_t    br_type,
    output logic        is_jump_op,

    output logic        is_imm,
    output logic [31:0] imm_b,
    output logic [31:0] imm_i,
    output logic [31:0] imm_s,
    output logic [31:0] imm_u,
    output logic [31:0] imm_j
);
    
    logic [4:0]  op;
    logic [2:0]  funct3;
    logic [6:0]  funct7;

    assign op = instr[6:2];
    assign is_imm = ~op[3];
    assign funct3 = instr[14:12];
    assign funct7 = instr[31:25];

    assign rd = instr[7+:4];
    assign rs1 = instr[15+:4];
    assign rs2 = instr[20+:4];

    // alu decode
    always_comb begin
        casez ({op,funct3})
            8'b00101_???,
            8'b0?000_???,
            8'b0?100_000 : alu_op = ADDER_OP;
            8'b0?100_010,
            8'b0?100_011,
            8'b11000_??? : alu_op = COMP_OP;
            8'b0?100_100 : alu_op = XOR_OP;
            8'b0?100_110 : alu_op = OR_OP;
            8'b0?100_111 : alu_op = AND_OP;
            8'b0?100_001,
            8'b0?100_101 : alu_op = SHIFTER_OP;
            default      : alu_op = ADDER_OP;
        endcase
    end

    // subtract enable
    always_comb begin
        casez ({op,funct3,funct7[5]})
            9'b01100_000_1,
            9'b0?100_010_?,
            9'b0?100_011_?,
            9'b11000_???_? : subtract = 1'b1;
            default        : subtract = 1'b0;
        endcase
    end

    assign is_auipc = (op == 5'b00101);

    // compare type decode
    assign comp_op = comp_t'(funct3);

    // shift type decode
    assign shift_right = funct3[2];
    assign shift_arith = funct7[5];

    // branch decode
    assign is_br_type = ({op[4:2]} == 3'b110);
    assign br_type = br_type_t'(op[3:2]);
    assign is_jump_op = is_br_type & op[0];

    // load/store decode
    assign is_load_op = (op == 5'b00000);
    assign load_op = load_op_t'(funct3);
    assign is_store_op = (op == 5'b01000);
    assign store_op = store_op_t'(funct3);

    // B-type: imm[12], imm[10:5], imm[4:1], imm[11] sign extended
    assign imm_b = {{19{instr[31]}}, instr[31], instr[7], instr[30:25], instr[11:8], 1'b0};
    // I-type: imm[11:0] sign extended
    assign imm_i = {{20{instr[31]}}, instr[31:20]};
    // S-type: imm[15:5] imm[4:0] sign extended
    assign imm_s = {{20{instr[31]}}, instr[31:25], instr[11:7]};
    // U-type: imm[31:12] lower 12 bits zero
    assign imm_u = {instr[31:12], 12'b0};
    // J-type: imm[20], imm[10:1], imm[11], imm[19:12]
    assign imm_j = {{11{instr[31]}}, instr[31], instr[19:12], instr[20], instr[30:21], 1'b0};

endmodule : decode
