module adder (
    input logic a,
    input logic a,
    output logic sum
);

    assign sum = a + b;

endmodule
