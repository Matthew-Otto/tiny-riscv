/home/ecelrc/students/cc75925/tiny-riscv/baseline/apr_run1/gscl45nm.lef